//: version "2.1-a1"
//: property encoding = "iso8859-1"
//: property locale = "en"
//: property prefix = "_GG"
//: property title = "rtm.v"
//: property timingViolationMode = 2
//: property initTime = "0 ns"

`timescale 1ns/1ns

//: /netlistBegin main
module main;    //: root_module
supply1 w7;    //: /sn:0 {0}(520,160)(520,121){1}
reg [3:0] w0;    //: /sn:0 {0}(#:107,68)(107,218)(234,218){1}
reg w29;    //: /sn:0 {0}(1092,58)(1103,58)(1103,127)(1044,127)(1044,192){1}
//: {2}(1046,194)(1155,194)(1155,215){3}
//: {4}(1044,196)(1044,314){5}
//: {6}(1046,316)(1159,316)(1159,340){7}
//: {8}(1044,318)(1044,760){9}
reg w30;    //: /sn:0 {0}(1221,760)(1221,259){1}
//: {2}(1223,257)(1268,257)(1268,273){3}
//: {4}(1221,255)(1221,130)(1177,130)(1177,111)(1044,111)(1044,58)(1036,58){5}
reg w12;    //: /sn:0 {0}(675,58)(693,58)(693,58)(692,58){1}
reg w10;    //: /sn:0 {0}(451,59)(465,59)(465,179)(483,179){1}
reg w31;    //: /sn:0 {0}(1238,59)(1248,59)(1248,145)(1096,145)(1096,444){1}
//: {2}(1098,446)(1162,446)(1162,471){3}
//: {4}(1096,448)(1096,608){5}
//: {6}(1098,610)(1162,610)(1162,633){7}
//: {8}(1096,612)(1096,760){9}
reg w33;    //: /sn:0 {0}(1182,59)(1190,59)(1190,120)(1237,120)(1237,522){1}
//: {2}(1239,524)(1268,524)(1268,543){3}
//: {4}(1237,526)(1237,760){5}
reg w14;    //: /sn:0 {0}(1408,57)(1431,57)(1431,317){1}
//: {2}(1429,319)(1382,319)(1382,374){3}
//: {4}(1431,321)(1431,356){5}
reg w11;    //: /sn:0 {0}(789,734)(789,741)(825,741)(825,585){1}
//: {2}(825,581)(825,433){3}
//: {4}(825,429)(825,280){5}
//: {6}(825,276)(825,132){7}
//: {8}(823,278)(789,278)(789,266){9}
//: {10}(823,431)(789,431)(789,421){11}
//: {12}(823,583)(789,583)(789,577){13}
reg w5;    //: /sn:0 {0}(203,58)(250,58)(250,205){1}
reg w9;    //: /sn:0 {0}(393,57)(401,57)(401,189)(483,189){1}
wire [3:0] w13;    //: /sn:0 {0}(#:1281,566)(1317,566)(1317,566)(1348,566){1}
//: {2}(1350,564)(1350,409){3}
//: {4}(1352,407)(1366,407){5}
//: {6}(1350,405)(1350,388){7}
//: {8}(1352,386)(#:1362,386)(1362,387)(1366,387){9}
//: {10}(1350,384)(#:1350,135){11}
//: {12}(1350,568)(1350,760){13}
wire w16;    //: /sn:0 {0}(655,766)(655,313){1}
//: {2}(657,311)(794,311)(794,345){3}
//: {4}(655,309)(655,180){5}
//: {6}(655,176)(655,135){7}
//: {8}(653,178)(536,178){9}
wire [3:0] w6;    //: /sn:0 {0}(1252,306)(1188,306)(1188,363)(#:1172,363){1}
wire w25;    //: /sn:0 {0}(784,345)(784,326)(753,326){1}
//: {2}(751,324)(751,172){3}
//: {4}(753,170)(784,170)(784,190){5}
//: {6}(751,168)(751,58)(708,58){7}
//: {8}(751,328)(751,485){9}
//: {10}(753,487)(784,487)(784,501){11}
//: {12}(751,489)(751,649)(784,649)(784,658){13}
wire [3:0] w4;    //: /sn:0 {0}(#:778,383)(311,383){1}
//: {2}(309,381)(#:309,230){3}
//: {4}(311,228)(778,228){5}
//: {6}(309,226)(309,177)(309,177)(309,135){7}
//: {8}(307,228)(#:263,228){9}
//: {10}(#:309,385)(309,537){11}
//: {12}(311,539)(778,539){13}
//: {14}(#:309,541)(309,694){15}
//: {16}(311,696)(778,696){17}
//: {18}(309,698)(309,753){19}
wire w36;    //: /sn:0 {0}(1472,135)(1472,419){1}
//: {2}(1470,421)(1431,421)(1431,404){3}
//: {4}(1472,423)(1472,758){5}
wire [3:0] w3;    //: /sn:0 {0}(1252,286)(1187,286)(1187,238)(#:1168,238){1}
wire [3:0] w20;    //: /sn:0 {0}(#:1307,135)(1307,213)(1307,213)(1307,294){1}
//: {2}(1305,296)(1295,296)(1295,296)(#:1281,296){3}
//: {4}(#:1307,298)(1307,362){5}
//: {6}(1309,364)(1417,364){7}
//: {8}(1307,366)(1307,758){9}
wire [3:0] w37;    //: /sn:0 {0}(#:1146,504)(940,504){1}
//: {2}(938,502)(938,385){3}
//: {4}(938,381)(938,250){5}
//: {6}(940,248)(1139,248){7}
//: {8}(938,246)(938,190)(938,190)(#:938,135){9}
//: {10}(936,383)(#:799,383){11}
//: {12}(938,506)(938,757){13}
wire w18;    //: /sn:0 {0}(794,658)(794,627)(717,627){1}
//: {2}(715,625)(715,204){3}
//: {4}(715,200)(715,135){5}
//: {6}(713,202)(536,202){7}
//: {8}(715,629)(715,767){9}
wire [3:0] w23;    //: /sn:0 {0}(1252,576)(1190,576)(1190,656)(#:1175,656){1}
wire [3:0] w21;    //: /sn:0 {0}(1252,556)(1189,556)(1189,494)(#:1175,494){1}
wire [3:0] w1;    //: /sn:0 {0}(#:799,696)(994,696){1}
//: {2}(996,694)(996,668){3}
//: {4}(998,666)(1146,666){5}
//: {6}(996,664)(996,375){7}
//: {8}(#:998,373)(1143,373){9}
//: {10}(996,371)(996,252)(996,252)(996,135){11}
//: {12}(996,698)(996,758){13}
wire [3:0] w32;    //: /sn:0 {0}(#:909,758)(909,486){1}
//: {2}(911,484)(#:1146,484){3}
//: {4}(909,482)(909,230){5}
//: {6}(911,228)(1139,228){7}
//: {8}(909,226)(909,180)(909,180)(#:909,135){9}
//: {10}(907,228)(#:799,228){11}
wire w8;    //: /sn:0 {0}(626,765)(626,168){1}
//: {2}(626,164)(626,154){3}
//: {4}(628,152)(794,152)(794,190){5}
//: {6}(626,150)(626,135){7}
//: {8}(624,166)(536,166){9}
wire w17;    //: /sn:0 {0}(684,766)(684,471){1}
//: {2}(686,469)(794,469)(794,501){3}
//: {4}(684,467)(684,192){5}
//: {6}(684,188)(684,135){7}
//: {8}(682,190)(536,190){9}
wire [3:0] w28;    //: /sn:0 {0}(#:1395,396)(1417,396){1}
wire [3:0] w2;    //: /sn:0 {0}(#:1446,380)(1522,380){1}
//: {2}(1524,378)(1524,255)(1524,255)(1524,135){3}
//: {4}(#:1524,382)(1524,776)(107,776)(107,238)(234,238){5}
wire [3:0] w15;    //: /sn:0 {0}(#:1146,646)(969,646){1}
//: {2}(967,644)(967,541){3}
//: {4}(967,537)(967,355){5}
//: {6}(969,353)(1143,353){7}
//: {8}(967,351)(967,242)(967,242)(#:967,135){9}
//: {10}(965,539)(#:799,539){11}
//: {12}(967,648)(967,758){13}
wire [1:0] w38;    //: /sn:0 {0}(#:489,184)(#:507,184){1}
//: enddecls

  //: LED clk3 (w18) @(715,128) /w:[ 5 ] /type:0
  //: joint g44 (w20) @(1307, 296) /w:[ -1 1 2 4 ]
  //: joint g8 (w18) @(715, 202) /w:[ -1 4 6 3 ]
  //: joint g4 (w2) @(1524, 380) /w:[ -1 2 1 4 ]
  //: VDD g16 (w7) @(531,121) /sn:0 /w:[ 1 ]
  //: joint g47 (w29) @(1044, 316) /w:[ 6 5 -1 8 ]
  //: joint g3 (w8) @(626, 166) /w:[ -1 2 8 1 ]
  //: joint g17 (w11) @(825, 583) /w:[ -1 2 12 1 ]
  //: joint g26 (w1) @(996, 696) /w:[ -1 2 1 12 ]
  //: SWITCH ctl_add (w5) @(186,58) /w:[ 0 ] /st:0 /dn:0
  _GGNDECODER4 #(4, 4) g2 (.I(w38), .E(w7), .Z0(w8), .Z1(w16), .Z2(w17), .Z3(w18));   //: @(520,184) /sn:0 /R:1 /w:[ 1 0 9 9 9 7 ] /ss:1 /do:1
  //: joint g30 (w4) @(309, 539) /w:[ 12 11 -1 14 ]
  //: joint g23 (w1) @(996, 373) /w:[ 8 10 -1 7 ]
  //: joint g24 (w15) @(967, 646) /w:[ 1 2 -1 12 ]
  //: joint g39 (w15) @(967, 539) /w:[ -1 4 10 3 ]
  //: SWITCH ctl_sa0 (w30) @(1019,58) /w:[ 5 ] /st:1 /dn:0
  _GGREG4 #(10, 10, 20) g1 (.Q(w32), .D(w4), .EN(w8), .CLR(w25), .CK(w11));   //: @(789,228) /sn:0 /R:1 /w:[ 11 5 5 5 9 ]
  //: joint g60 (w14) @(1431, 319) /w:[ -1 1 2 4 ]
  //: SWITCH ctl_sb1 (w31) @(1221,59) /w:[ 0 ] /st:1 /dn:0
  //: joint g29 (w4) @(309, 383) /w:[ 1 2 -1 10 ]
  //: LED reg0 (w32) @(909,128) /w:[ 9 ] /type:2
  //: LED reg2 (w15) @(967,128) /w:[ 9 ] /type:2
  //: SWITCH ctl_clear (w12) @(658,58) /w:[ 0 ] /st:0 /dn:0
  //: LED g51 (w2) @(1524,128) /sn:0 /w:[ 3 ] /type:2
  //: joint g18 (w11) @(825, 431) /w:[ -1 4 10 3 ]
  //: LED reg3 (w1) @(996,128) /w:[ 11 ] /type:2
  //: LED carry_out (w36) @(1472,128) /w:[ 0 ] /type:0
  //: joint g25 (w37) @(938, 383) /w:[ -1 4 10 3 ]
  _GGREG4 #(10, 10, 20) g10 (.Q(w37), .D(w4), .EN(w16), .CLR(w25), .CK(w11));   //: @(789,383) /sn:0 /R:1 /w:[ 11 0 3 0 11 ]
  //: LED clk1 (w16) @(655,128) /w:[ 7 ] /type:0
  //: LED clk2 (w17) @(684,128) /w:[ 7 ] /type:0
  //: joint g49 (w30) @(1221, 257) /w:[ 2 4 -1 1 ]
  //: joint g6 (w16) @(655, 178) /w:[ -1 6 8 5 ]
  //: joint g50 (w33) @(1237, 524) /w:[ 2 1 -1 4 ]
  //: LED reg1 (w37) @(938,128) /w:[ 9 ] /type:2
  //: joint g58 (w18) @(715, 627) /w:[ 1 2 -1 8 ]
  //: joint g56 (w17) @(684, 469) /w:[ 2 4 -1 1 ]
  _GGMUX2x4 #(8, 8) g35 (.I0(w32), .I1(w37), .S(w31), .Z(w21));   //: @(1162,494) /sn:0 /R:1 /w:[ 3 0 3 1 ] /ss:1 /do:1
  //: joint g7 (w17) @(684, 190) /w:[ -1 6 8 5 ]
  //: joint g9 (w32) @(909, 228) /w:[ 6 8 10 5 ]
  //: joint g59 (w13) @(1350, 407) /w:[ 4 6 -1 3 ]
  //: joint g22 (w37) @(938, 504) /w:[ 1 2 -1 12 ]
  _GGMUX2x4 #(8, 8) g31 (.I0(w3), .I1(w6), .S(w30), .Z(w20));   //: @(1268,296) /sn:0 /R:1 /w:[ 0 0 3 3 ] /ss:1 /do:1
  _GGMUX2x4 #(8, 10) g45 (.I0(w13), .I1(~w13), .S(w14), .Z(w28));   //: @(1382,397) /sn:0 /R:1 /w:[ 5 9 3 0 ] /ss:1 /do:0
  //: joint g54 (w8) @(626, 152) /w:[ 4 6 -1 3 ]
  _GGMUX2x4 #(8, 8) g33 (.I0(w32), .I1(w37), .S(w29), .Z(w3));   //: @(1155,238) /sn:0 /R:1 /w:[ 7 7 3 1 ] /ss:1 /do:1
  //: joint g41 (w13) @(1350, 566) /w:[ -1 2 1 12 ]
  _GGMUX2x4 #(8, 8) g36 (.I0(w15), .I1(w1), .S(w31), .Z(w23));   //: @(1162,656) /sn:0 /R:1 /w:[ 0 5 7 1 ] /ss:1 /do:1
  //: LED a_bus (w20) @(1307,128) /w:[ 0 ] /type:2
  //: LED clk0 (w8) @(626,128) /w:[ 7 ] /type:0
  //: joint g40 (w1) @(996, 666) /w:[ 4 6 -1 3 ]
  //: joint g42 (w20) @(1307, 364) /w:[ 6 5 -1 8 ]
  assign w38 = {w9, w10}; //: CONCAT g52  @(488,184) /sn:0 /w:[ 0 1 1 ] /dr:1 /tp:0 /drp:1
  _GGREG4 #(10, 10, 20) g12 (.Q(w1), .D(w4), .EN(w18), .CLR(w25), .CK(w11));   //: @(789,696) /sn:0 /R:1 /w:[ 0 17 0 13 0 ]
  //: SWITCH ctl_sa1 (w29) @(1075,58) /w:[ 0 ] /st:0 /dn:0
  //: DIP indata (w0) @(107,58) /w:[ 0 ] /st:2 /dn:0
  //: joint g46 (w4) @(309, 696) /w:[ 16 15 -1 18 ]
  //: SWITCH carry_in (w14) @(1391,57) /w:[ 0 ] /st:1 /dn:0
  //: joint g57 (w36) @(1472, 421) /w:[ -1 1 2 4 ]
  //: joint g28 (w4) @(309, 228) /w:[ 4 6 8 3 ]
  _GGMUX2x4 #(8, 8) g34 (.I0(w15), .I1(w1), .S(w29), .Z(w6));   //: @(1159,363) /sn:0 /R:1 /w:[ 7 9 7 1 ] /ss:1 /do:1
  //: joint g5 (w11) @(825, 278) /w:[ -1 6 8 5 ]
  //: joint g14 (w25) @(751, 326) /w:[ 1 2 -1 8 ]
  //: SWITCH ctl_d0 (w9) @(376,57) /w:[ 0 ] /st:1 /dn:0
  _GGREG4 #(10, 10, 20) g11 (.Q(w15), .D(w4), .EN(w17), .CLR(w25), .CK(w11));   //: @(789,539) /sn:0 /R:1 /w:[ 11 13 3 11 13 ]
  //: SWITCH ctl_d1 (w10) @(434,59) /w:[ 0 ] /st:1 /dn:0
  //: joint g21 (w15) @(967, 353) /w:[ 6 8 -1 5 ]
  //: LED b_bus (w13) @(1350,128) /w:[ 11 ] /type:2
  //: joint g19 (w37) @(938, 248) /w:[ 6 8 -1 5 ]
  //: joint g20 (w32) @(909, 484) /w:[ 2 4 -1 1 ]
  _GGMUX2x4 #(8, 8) g32 (.I0(w21), .I1(w23), .S(w33), .Z(w13));   //: @(1268,566) /sn:0 /R:1 /w:[ 0 0 3 0 ] /ss:1 /do:1
  _GGMUX2x4 #(8, 8) g0 (.I0(w0), .I1(w2), .S(w5), .Z(w4));   //: @(250,228) /sn:0 /R:1 /w:[ 1 5 1 9 ] /ss:1 /do:1
  _GGADD4 #(36, 38, 30, 32) g43 (.A(w28), .B(w20), .S(w2), .CI(w14), .CO(w36));   //: @(1433,380) /sn:0 /R:1 /w:[ 1 7 0 5 3 ]
  //: SWITCH ctl_sb0 (w33) @(1165,59) /w:[ 0 ] /st:1 /dn:0
  //: joint g15 (w25) @(751, 487) /w:[ 10 9 -1 12 ]
  //: joint g38 (w31) @(1096, 446) /w:[ 2 1 -1 4 ]
  //: joint g48 (w31) @(1096, 610) /w:[ 6 5 -1 8 ]
  _GGNBUF #(2) g27 (.I(w12), .Z(w25));   //: @(698,58) /sn:0 /w:[ 1 7 ]
  //: LED d_bus (w4) @(309,128) /w:[ 7 ] /type:2
  //: joint g37 (w29) @(1044, 194) /w:[ 2 1 -1 4 ]
  //: joint g55 (w16) @(655, 311) /w:[ 2 4 -1 1 ]
  //: joint g53 (w13) @(1350, 386) /w:[ 8 10 -1 7 ]
  //: SWITCH clock (w11) @(825,119) /R:3 /w:[ 7 ] /st:0 /dn:0
  //: joint g13 (w25) @(751, 170) /w:[ 4 6 -1 3 ]

endmodule
//: /netlistEnd

